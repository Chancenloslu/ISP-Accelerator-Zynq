package Settings;
//  Integer width = 1173;
//  Integer height = 470;
  Integer width = 260;
  Integer height = 260;
  Integer n_vals = width * height;
  Integer n_out = (width-2) * (height-2);

typedef 32 F_AW;
typedef 128 F_RD_DW;
typedef 128 F_WR_DW;
typedef 2 F_ID_W;
typedef 2 F_USER_W;
  
typedef 5 L_AW;
typedef 32 L_DW;

endpackage
