package MyTypes;
import Vector :: *;
typedef Bit#(8) GrayScale;
typedef Bit#(24) RGB;
typedef Vector#(3, Bit#(8)) Field_RGB;

endpackage
